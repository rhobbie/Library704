// Verilog test bench for SYSTEM
`timescale 100ns/100ns
module SYSTEM_tb;

reg CL=0;
reg RESET=1;

SYSTEM S(CL,RESET);

integer i;

initial 
begin
  
  $dumpfile("Sort.vcd");
  $dumpvars(0, SYSTEM_tb);   
  
  # 5 RESET=0;
  for(i=0;i<12000;i=i+1)
  begin
    # 5 CL=1;
    # 5 CL=0;   
  end
  
end

initial
begin  
  # 10000
  
S.SP.Mem['o00000]=36'o0_53400_2_00015; //         LXA CONST,2      Set count of no. of passes
S.SP.Mem['o00001]=36'o4_53400_1_00010; //  PASS   LXD SKIP,1       Consider 1st pair
S.SP.Mem['o00002]=36'o4_63400_2_00011; //         SXD TEST,2       Set test for end of pass.
S.SP.Mem['o00003]=36'o0_56000_1_00016; //  NEXT   LDQ A,1
S.SP.Mem['o00004]=36'o0_50000_1_00017; //         CLA A+1,1
S.SP.Mem['o00005]=36'o0_04000_0_00010; //         TLQ SKIP         is the pair out-of-order?
S.SP.Mem['o00006]=36'o0_60100_1_00016; //         STO A,1          yes, interchange them
S.SP.Mem['o00007]=36'o4_60000_1_00017; //         STQ A+1,1
S.SP.Mem['o00010]=36'o1_77777_1_00011; //  SKIP   TXI SKIP+1,1,-1  Consider next pair
S.SP.Mem['o00011]=36'o3_00000_1_00003; //  TEST   TXH NEXT,1,-     go NEXT if not end
S.SP.Mem['o00012]=36'o1_00001_2_00013; //  Q      TXI Q+1,2,1      Prepare for next pass
S.SP.Mem['o00013]=36'o7_77776_2_00001; //         TXL PASS,2,-2    Go beck for next pass, or
S.SP.Mem['o00014]=36'o0_42000_0_00000; //         HPR              stop
S.SP.Mem['o00015]=36'o0_00000_0_77766; //  CONST  PZE -10          Adress has 2^15-10=32758
S.SP.Mem['o00016]=36'o0_00000_0_00010; //  A      PZE 0
S.SP.Mem['o00017]=36'o0_00000_0_00004; //         PZE 4
S.SP.Mem['o00020]=36'o0_00000_0_11471; //         PZE 4921
S.SP.Mem['o00021]=36'o0_00000_0_00042; //         PZE 34
S.SP.Mem['o00022]=36'o0_00000_0_04662; //         PZE 2482
S.SP.Mem['o00023]=36'o0_00000_0_00501; //         PZE 321
S.SP.Mem['o00024]=36'o0_00000_0_04436; //         PZE 2334
S.SP.Mem['o00025]=36'o0_00000_0_00143; //         PZE 99
S.SP.Mem['o00026]=36'o0_00000_0_04243; //         PZE 2211
S.SP.Mem['o00027]=36'o0_00000_0_00173; //         PZE 123
S.SP.Mem['o00030]=36'o0_00000_0_00301; //         PZE 193
  
  #  1000  
      S.OP.START_BUTTON.State=1;
  # 10000  
      S.OP.START_BUTTON.State=0;  
   # 120000      
    ;

end
wire [35:0] A1,A2,A3,A4,A5,A6,A7,A8,A9,A10;
assign A1=S.SP.Mem['o00017];
assign A2=S.SP.Mem['o00020];
assign A3=S.SP.Mem['o00021];
assign A4=S.SP.Mem['o00022];
assign A5=S.SP.Mem['o00023];
assign A6=S.SP.Mem['o00024];
assign A7=S.SP.Mem['o00025];
assign A8=S.SP.Mem['o00026];
assign A9=S.SP.Mem['o00027];
assign A10=S.SP.Mem['o00030];


wire PROG_STOP;
assign PROG_STOP=S.OP.PROG_STOP_LITE.State;

wire  ACC_OVERFLOW;
assign ACC_OVERFLOW=S.OP.ACC_OVERFLOW_LITE.State;

wire DIV_CHECK;
assign DIV_CHECK=S.OP.DIV_CHECK.State;

wire RD_WR_SELECT;
assign RD_WR_SELECT=S.OP.RD_WR_SELECT.State;

wire MQ_OV;
assign MQ_OV=S.OP.MQ_OV_LITE.State;

wire RD_WR_CHECK;
assign RD_WR_CHECK=S.OP.RD_WR_CHECK.State;


wire [12:0] XR;

assign XR={S.OP.XR_COL_0_NEON.State,S.OP.XR_COL_1_NEON.State,S.OP.XR_COL_2_NEON.State,S.OP.XR_COL_3_NEON.State,S.OP.XR_COL_4_NEON.State,S.OP.XR_COL_5_NEON.State,
  S.OP.XR_COL_6_NEON.State,S.OP.XR_COL_7_NEON.State,S.OP.XR_COL_8_NEON.State,S.OP.XR_COL_9_NEON.State,S.OP.XR_COL_10_NEON.State,S.OP.XR_COL_11_NEON.State,     
  S.OP.XR_COL_12_NEON.State};

wire TAPE_CHECK;
assign TAPE_CHECK=S.OP.TAPE_CHECK_NEON.State;


wire READY;
assign READY=S.OP.READY_LIGHT.State;

wire AUTO;
assign AUTO=S.OP.AUTO_LIGHT.State;


wire  [35:0] STG;
assign STG={S.OP.STG_S_NEON.State,S.OP.STG_1_NEON.State,S.OP.STG_2_NEON.State,S.OP.STG_3_NEON.State,S.OP.STG_4_NEON.State,S.OP.STG_5_NEON.State,
  S.OP.STG_6_NEON.State,S.OP.STG_7_NEON.State,S.OP.STG_8_NEON.State,S.OP.STG_9_NEON.State,S.OP.STG_10_NEON.State,S.OP.STG_11_NEON.State,     
  S.OP.STG_12_NEON.State,S.OP.STG_13_NEON.State,S.OP.STG_14_NEON.State,S.OP.STG_15_NEON.State,S.OP.STG_16_NEON.State,S.OP.STG_17_NEON.State,
  S.OP.STG_18_NEON.State,S.OP.STG_19_NEON.State,S.OP.STG_20_NEON.State,S.OP.STG_21_NEON.State,S.OP.STG_22_NEON.State,S.OP.STG_23_NEON.State,
  S.OP.STG_24_NEON.State,S.OP.STG_25_NEON.State,S.OP.STG_26_NEON.State,S.OP.STG_27_NEON.State,S.OP.STG_28_NEON.State,S.OP.STG_29_NEON.State,
  S.OP.STG_30_NEON.State,S.OP.STG_31_NEON.State,S.OP.STG_32_NEON.State,S.OP.STG_33_NEON.State,S.OP.STG_34_NEON.State,S.OP.STG_35_NEON.State};


wire  [37:0] ACC;
assign ACC={S.OP.ACC_S_NEON.State,S.OP.ACC_Q_NEON.State,S.OP.ACC_P_NEON.State,S.OP.ACC_1_NEON.State,S.OP.ACC_2_NEON.State,S.OP.ACC_3_NEON.State,S.OP.ACC_4_NEON.State,S.OP.ACC_5_NEON.State,
  S.OP.ACC_6_NEON.State,S.OP.ACC_7_NEON.State,S.OP.ACC_8_NEON.State,S.OP.ACC_9_NEON.State,S.OP.ACC_10_NEON.State,S.OP.ACC_11_NEON.State,     
  S.OP.ACC_12_NEON.State,S.OP.ACC_13_NEON.State,S.OP.ACC_14_NEON.State,S.OP.ACC_15_NEON.State,S.OP.ACC_16_NEON.State,S.OP.ACC_17_NEON.State,
  S.OP.ACC_18_NEON.State,S.OP.ACC_19_NEON.State,S.OP.ACC_20_NEON.State,S.OP.ACC_21_NEON.State,S.OP.ACC_22_NEON.State,S.OP.ACC_23_NEON.State,
  S.OP.ACC_24_NEON.State,S.OP.ACC_25_NEON.State,S.OP.ACC_26_NEON.State,S.OP.ACC_27_NEON.State,S.OP.ACC_28_NEON.State,S.OP.ACC_29_NEON.State,
  S.OP.ACC_30_NEON.State,S.OP.ACC_31_NEON.State,S.OP.ACC_32_NEON.State,S.OP.ACC_33_NEON.State,S.OP.ACC_34_NEON.State,S.OP.ACC_35_NEON.State};

wire  [35:0] MQ;
assign MQ={S.OP.MQ_S_NEON.State,S.OP.MQ_1_NEON.State,S.OP.MQ_2_NEON.State,S.OP.MQ_3_NEON.State,S.OP.MQ_4_NEON.State,S.OP.MQ_5_NEON.State,
  S.OP.MQ_6_NEON.State,S.OP.MQ_7_NEON.State,S.OP.MQ_8_NEON.State,S.OP.MQ_9_NEON.State,S.OP.MQ_10_NEON.State,S.OP.MQ_11_NEON.State,     
  S.OP.MQ_12_NEON.State,S.OP.MQ_13_NEON.State,S.OP.MQ_14_NEON.State,S.OP.MQ_15_NEON.State,S.OP.MQ_16_NEON.State,S.OP.MQ_17_NEON.State,
  S.OP.MQ_18_NEON.State,S.OP.MQ_19_NEON.State,S.OP.MQ_20_NEON.State,S.OP.MQ_21_NEON.State,S.OP.MQ_22_NEON.State,S.OP.MQ_23_NEON.State,
  S.OP.MQ_24_NEON.State,S.OP.MQ_25_NEON.State,S.OP.MQ_26_NEON.State,S.OP.MQ_27_NEON.State,S.OP.MQ_28_NEON.State,S.OP.MQ_29_NEON.State,
  S.OP.MQ_30_NEON.State,S.OP.MQ_31_NEON.State,S.OP.MQ_32_NEON.State,S.OP.MQ_33_NEON.State,S.OP.MQ_34_NEON.State,S.OP.MQ_35_NEON.State};


wire  [12:0] INST_CTR;
assign INST_CTR={S.OP.INST_CTR_5_NEON.State,
 S.OP.INST_CTR_6_NEON.State,S.OP.INST_CTR_7_NEON.State,S.OP.INST_CTR_8_NEON.State,S.OP.INST_CTR_9_NEON.State,S.OP.INST_CTR_10_NEON.State,S.OP.INST_CTR_11_NEON.State,
 S.OP.INST_CTR_12_NEON.State,S.OP.INST_CTR_13_NEON.State,S.OP.INST_CTR_14_NEON.State,S.OP.INST_CTR_15_NEON.State,S.OP.INST_CTR_16_NEON.State,S.OP.INST_CTR_17_NEON.State};  

wire TRAP_MODE;
assign TRAP_MODE=S.OP.TRAP_MODE_NEON.State;

 
wire  [17:0] INST_REG;
assign INST_REG={S.OP.INST_REG_S_NEON.State,S.OP.INST_REG_1_NEON.State,S.OP.INST_REG_2_NEON.State,S.OP.INST_REG_3_NEON.State,S.OP.INST_REG_4_NEON.State,S.OP.INST_REG_5_NEON.State,
  S.OP.INST_REG_6_NEON.State,S.OP.INST_REG_7_NEON.State,S.OP.INST_REG_8_NEON.State,S.OP.INST_REG_9_NEON.State,S.OP.INST_REG_10_NEON.State,S.OP.INST_REG_11_NEON.State,     
  S.OP.INST_REG_12_NEON.State,S.OP.INST_REG_13_NEON.State,S.OP.INST_REG_14_NEON.State,S.OP.INST_REG_15_NEON.State,S.OP.INST_REG_16_NEON.State,S.OP.INST_REG_17_NEON.State};

wire SENSE_LIGHT_1;
assign SENSE_LIGHT_1=S.OP.SENSE_LIGHT_1_NEON.State;

wire SENSE_LIGHT_2;
assign SENSE_LIGHT_2=S.OP.SENSE_LIGHT_2_NEON.State;

wire SENSE_LIGHT_3;
assign SENSE_LIGHT_3=S.OP.SENSE_LIGHT_3_NEON.State;

wire SENSE_LIGHT_4;
assign SENSE_LIGHT_4=S.OP.SENSE_LIGHT_4_NEON.State;

wire [12:0] XRA;
wire [12:0] XRB;
wire [12:0] XRC;
assign XRA={S.MF4.A36._03O,S.MF4.A07_7,S.MF4.A08_7,S.MF4.A09_7,S.MF4.C07_7,S.MF4.C08_7,S.MF4.C09_7,S.MF4.D07_7,S.MF4.D08_7,S.MF4.D09_7,S.MF4.E07_7,S.MF4.E08_7,S.MF4.E09_7};
assign XRB={S.MF4.A36._04O,S.MF4.A10_7,S.MF4.A11_7,S.MF4.A13_7,S.MF4.C10_7,S.MF4.C11_7,S.MF4.C13_7,S.MF4.D10_7,S.MF4.D11_7,S.MF4.D13_7,S.MF4.E10_7,S.MF4.E11_7,S.MF4.E13_7};
assign XRC={S.MF4.A36._06O,S.MF4.A14_7,S.MF4.A15_7,S.MF4.A16_7,S.MF4.C14_7,S.MF4.C15_7,S.MF4.C16_7,S.MF4.D14_7,S.MF4.D15_7,S.MF4.D16_7,S.MF4.E14_7,S.MF4.E15_7,S.MF4.E16_7};

wire [37:0] adder_input;

assign adder_input={S.MF2.D01_7,S.MF2.D02_7,S.MF2.A04._04BO,S.MF2.A05._04BO,S.MF2.A06._04BO,S.MF2.A07._04BO,S.MF2.A08._04BO,S.MF2.A09._04BO,S.MF2.A10._04BO,S.MF2.A11._04BO,S.MF2.A12._04BO,
S.MF2.A13._04BO,S.MF2.A14._04BO,S.MF2.A15._04BO,S.MF2.A16._04BO,S.MF2.A17._04BO,S.MF2.A18._04BO,S.MF2.A19._04BO,S.MF2.A20._04BO,S.MF2.A21._04BO,S.MF2.A22._04BO,S.MF2.A23._04BO,
S.MF2.A24._04BO,S.MF2.A25._04BO,S.MF2.A26._04BO,S.MF2.A27._04BO,S.MF2.A28._04BO,S.MF2.A29._04BO,S.MF2.A30._04BO,S.MF2.A31._04BO,S.MF2.A32._04BO,S.MF2.A33._04BO,S.MF2.A34._04BO,
S.MF2.A35._04BO,S.MF2.A36._04BO,S.MF2.A37._04BO,S.MF2.A38._04BO};

wire [37:0] carry_in;

assign carry_in={S.MF2.C01_7,S.MF2.C02_7,S.MF2.B04_2,S.MF2.B05_2,S.MF2.B06_2,S.MF2.B07_2,S.MF2.B08_2,S.MF2.B09_2,S.MF2.B10_2,S.MF2.B11_2,S.MF2.B12_2,S.MF2.B13_2,S.MF2.B14_2,S.MF2.B15_2,
S.MF2.B16_2,S.MF2.B17_2,S.MF2.B18_7_i,S.MF2.B19_7_i,S.MF2.B20_2,S.MF2.B21_2,S.MF2.B22_2,S.MF2.B23_2,S.MF2.B24_2,S.MF2.B25_2,S.MF2.B26_2,S.MF2.B27_2,S.MF2.B28_2,S.MF2.B29_2,S.MF2.B30_2,
S.MF2.B31_2,S.MF2.B32_2,S.MF2.B33_2,S.MF2.B34_2,S.MF2.B35_2,S.MF2.B36_2,S.MF2.B37_2,S.MF2.B38_2};

wire [37:0] input_t_c;
assign input_t_c={S.MF2.A01._03AO,S.MF2.A02._03BO,S.MF2.A04._04AO,S.MF2.A05._04AO,S.MF2.A06._04AO,S.MF2.A07._04AO,S.MF2.A08._04AO,S.MF2.A09._04AO,S.MF2.A10._04AO,S.MF2.A11._04AO,
S.MF2.A12._04AO,S.MF2.A13._04AO,S.MF2.A14._04AO,S.MF2.A15._04AO,S.MF2.A16._04AO,S.MF2.A17._04AO,S.MF2.A18._04AO,S.MF2.A19._04AO,S.MF2.A20._04AO,S.MF2.A21._04AO,S.MF2.A22._04AO,
S.MF2.A23._04AO,S.MF2.A24._04AO,S.MF2.A25._04AO,S.MF2.A26._04AO,S.MF2.A27._04AO,S.MF2.A28._04AO,S.MF2.A29._04AO,S.MF2.A30._04AO,S.MF2.A31._04AO,S.MF2.A32._04AO,S.MF2.A33._04AO,
S.MF2.A34._04AO,S.MF2.A35._04AO,S.MF2.A36._04AO,S.MF2.A37._04AO,S.MF2.A38._04AO};

wire [37:0] carry_out;
assign carry_out={S.MF2.C01_2,S.MF2.C02_2,S.MF2.B04_6,S.MF2.B05_6,S.MF2.B06_6,S.MF2.B07_6,S.MF2.B08_6,S.MF2.B09_6,S.MF2.B10_6,S.MF2.B11_6,S.MF2.B12_6,S.MF2.B13_6,S.MF2.B14_6,S.MF2.B15_6,
S.MF2.B16_6,S.MF2.B17_6,S.MF2.B18_6,S.MF2.B19_6,S.MF2.B20_6,S.MF2.B21_6_o,S.MF2.B22_6,S.MF2.B23_6,S.MF2.B24_6,S.MF2.B25_6,S.MF2.B26_6,S.MF2.B27_6,S.MF2.B28_6,S.MF2.B29_6,S.MF2.B30_6,
S.MF2.B31_6,S.MF2.B32_6,S.MF2.B33_6,S.MF2.B34_6,S.MF2.B35_6,S.MF2.B36_6,S.MF2.B37_6,S.MF2.B38_6};

wire [37:0] sum_out;
assign sum_out={S.MF2.E01_3,S.MF2.D02_8,S.MF2.D04_8,S.MF2.D05_8,S.MF2.D06_8,S.MF2.D07_8,S.MF2.D08_8,S.MF2.D09_8,S.MF2.D10_8,S.MF2.D11_8,S.MF2.D12_8,S.MF2.D13_8,S.MF2.D14_8,S.MF2.D15_8,
S.MF2.D16_8,S.MF2.D17_8,S.MF2.D18_8,S.MF2.D19_8,S.MF2.D20_8,S.MF2.D21_8,S.MF2.D22_8,S.MF2.D23_8,S.MF2.D24_8,S.MF2.D25_8,S.MF2.D26_8,S.MF2.D27_8,S.MF2.D28_8,S.MF2.D29_8,S.MF2.D30_8,
S.MF2.D31_8,S.MF2.D32_8,S.MF2.D33_8,S.MF2.D34_8,S.MF2.D35_8,S.MF2.D36_8,S.MF2.D37_8,S.MF2.D38_8};

endmodule